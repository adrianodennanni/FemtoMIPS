-------------------------------------------------------------------------------
--
-- Title       : PROC
-- Design      : femtomips
-- Author      : adrianodennanni@hotmail.com
-- Company     : USP
--
-------------------------------------------------------------------------------
--
-- File        : C:\Users\adria\Desktop\FemtoMIPS\femtomips\compile\PROC.vhd
-- Generated   : Sun Jul  3 17:16:46 2016
-- From        : C:\Users\adria\Desktop\FemtoMIPS\femtomips\src\PROC.bde
-- By          : Bde2Vhdl ver. 2.6
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------
-- Design unit header --
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_signed.all;
use IEEE.std_logic_unsigned.all;


entity PROC is 
end PROC;

architecture PROC of PROC is

begin

end PROC;
