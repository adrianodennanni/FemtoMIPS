-------------------------------------------------------------------------------
--
-- Title       : No Title
-- Design      : Biblioteca_de_Componentes
-- Author      : LARC
-- Company     : LARC
--
-------------------------------------------------------------------------------
--
-- File        : c:\Arquivos de programas\Aldec\Active-HDL 8.2\Vlib\Biblioteca_de_Componentes\compile\#LARC.vhd
-- Generated   : Thu Aug 26 15:57:11 2010
-- From        : c:\Arquivos de programas\Aldec\Active-HDL 8.2\Vlib\Biblioteca_de_Componentes\src\#LARC.bde
-- By          : Bde2Vhdl ver. 2.6
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------
-- Design unit header --
library IEEE;
use IEEE.std_logic_1164.all;


entity \#LARC\ is 
end \#LARC\;

architecture \#LARC\ of \#LARC\ is

begin

end \#LARC\;
